//module tanh#(parameter width = 10)
//			  (value,
//			   clk,
//				tanh_val);