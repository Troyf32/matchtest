// megafunction wizard: %ALTSQRT%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTSQRT 

// ============================================================
// File Name: sqrt_16bit.v
// Megafunction Name(s):
// 			ALTSQRT
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 13.1.0 Build 162 10/23/2013 SJ Web Edition
// ************************************************************


//Copyright (C) 1991-2013 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module sqrt_16bit (
	clk,
	radical,
	q,
	remainder);

	input	  clk;
	input	[15:0]  radical;
	output	[7:0]  q;
	output	[8:0]  remainder;

	wire [7:0] sub_wire0;
	wire [8:0] sub_wire1;
	wire [7:0] q = sub_wire0[7:0];
	wire [8:0] remainder = sub_wire1[8:0];

	altsqrt	ALTSQRT_component (
				.clk (clk),
				.radical (radical),
				.q (sub_wire0),
				.remainder (sub_wire1)
				// synopsys translate_off
				,
				.aclr (),
				.ena ()
				// synopsys translate_on
				);
	defparam
		ALTSQRT_component.pipeline = 4,
		ALTSQRT_component.q_port_width = 8,
		ALTSQRT_component.r_port_width = 9,
		ALTSQRT_component.width = 16;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: PIPELINE NUMERIC "4"
// Retrieval info: CONSTANT: Q_PORT_WIDTH NUMERIC "8"
// Retrieval info: CONSTANT: R_PORT_WIDTH NUMERIC "9"
// Retrieval info: CONSTANT: WIDTH NUMERIC "16"
// Retrieval info: USED_PORT: clk 0 0 0 0 INPUT NODEFVAL "clk"
// Retrieval info: USED_PORT: q 0 0 8 0 OUTPUT NODEFVAL "q[7..0]"
// Retrieval info: USED_PORT: radical 0 0 16 0 INPUT NODEFVAL "radical[15..0]"
// Retrieval info: USED_PORT: remainder 0 0 9 0 OUTPUT NODEFVAL "remainder[8..0]"
// Retrieval info: CONNECT: @clk 0 0 0 0 clk 0 0 0 0
// Retrieval info: CONNECT: @radical 0 0 16 0 radical 0 0 16 0
// Retrieval info: CONNECT: q 0 0 8 0 @q 0 0 8 0
// Retrieval info: CONNECT: remainder 0 0 9 0 @remainder 0 0 9 0
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_16bit.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_16bit.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_16bit.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_16bit.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_16bit_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_16bit_bb.v FALSE
// Retrieval info: LIB_FILE: altera_mf
